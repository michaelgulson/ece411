//insert top level for mp3 here
import rv32i_types::*;

module mp3
(
    input rst,
    input pmem_resp,
    input [63:0] pmem_rdata,
    output logic pmem_read,
    output logic pmem_write,
    output rv32i_word pmem_address,
    output [63:0] pmem_wdata
);
cpu cpu(

);
cache i_cache(

); 
cache d_cache(

);
cache l2_cache(

);

endmodule : mp3