module PHT #(n)