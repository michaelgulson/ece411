//more caches to come