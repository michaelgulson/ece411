//insert top level for mp3 here